----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 19.02.2019 11:40:34
-- Design Name: 
-- Module Name: full_adder - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity full_adder is
    port (
        x, y, z : in std_logic;
        s, c : out std_logic
        );
end full_adder;

architecture Behavioral of full_adder is

    component half_adder
        port(
            x, y : in std_logic;
            s, c : out std_logic
            );
    end component;
    
    signal hs, hc, tc: std_logic;
    begin
        HA1: half_adder port map (
            x=>x, y=>y, s=>hs, c=>hc
        );
        HA2: half_adder port map (
             x=>hs, y=>z, s=>s, c=>tc
        );
        
        c <= tc or hc;
    


end Behavioral;
